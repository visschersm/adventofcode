module y2015

pub struct Solution01 {

}

pub fn (s Solution01) part1(input_file string) {
	println("Part1 not yet implemented")
}

pub fn (s Solution01) part2(input_file string) {
	println("Part2 not yet implemented")
}